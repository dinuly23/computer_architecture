// ******************************
// *модуль register_sload_sreset*
// ******************************
// = Входы =
// [шина] i   [W]: входные данные
// [бит ] l      : синхронный сигнал загрузки (сохранения входных данных по переднему фронту clk)
// [бит ] clk    : тактовый сигнал
// [бит ] rst    : синхронный сигнал сброса: сохранить значение по умолчанию по переднему фронту clk
//
// = Выходы =
// [шина] o [W]: выходные данные: непрерывно выводится последнее сохранённое значение
//
// = Параметры =
// W  [16]: ширина шин входных и выходных данных
// DV [ 0]: значение по умолчанию, сохраняемое при сбросе
//
// = Функционирование =
// В выходную шину непрерывно выводится последнее сохранённое значение.
// Значение сохраняется по каждому переднему фронту clk:
// * если "rst == 1", то сохраняется значение DV;
// * иначе сохраняется значение i.
// До первого переднего фронта сигнала clk сохранённое значение не определено (x).
module register_sload_sreset(i, l, clk, rst, o);
  parameter W = 16;
  parameter DV = 0;
  input [W-1:0] i;
  input l, clk, rst;
  output reg [W-1:0] o;
  
  always @(posedge clk)
    if(rst) o <= DV;
    else if(l) o <= i;
endmodule
