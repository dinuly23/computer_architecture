// ************
// *модуль mux*
// ************
// = Входы =
// [шина] i [DW*(2**CW)]: шина, разбитая на 2**CW блоков b(k) ширины DW: i = {b(0), b(1), ..., b(2**CW-1)}; ровно один из этих блоков перенаправляется на выход
// [шина] s [CW        ]: двоичная запись номера блока, перенаправляемого на выход
//
// = Выходы =
// [шина] o [DW]: непрерывно выводится значение блока b(s)
//
// = Параметры =
// DW [1]: ширина информационной шины o и блоков b(k)
// CW [2]: ширина управляющей шины s и логарифм количества блоков b(k)
module mux(i, s, o);
  parameter DW = 1;
  parameter CW = 2;
  localparam N = 2**CW;
  input [DW*N-1:0] i;
  input [CW-1:0] s;
  output [DW-1:0] o;
  
  wire [DW-1:0] b[0:N-1];
  
  genvar k;
  for(k = 0; k < N; k = k + 1)
    assign b[k] = i[DW*(N-k)-1:DW*(N-1-k)];
  
  assign o = b[s];
endmodule
