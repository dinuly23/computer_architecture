// **************
// *модуль demux*
// **************
// = Входы =
// [шина] i [DW]: значение этой шины непрерывно перенаправляется на выход
// [шина] s [CW]: двоичная запись номера блока выходной шины, в который надо перенаправить i
//
// = Выходы =
// [шина] o [DW*(2**CW)]:
//   * шина разбита на 2**CW блоков b(k) ширины DW: o = {b(0), b(1), ..., b(2**CW-1)}
//   * вход i непрерывно перенаправляется на блок b(s)
//   * в остальные блоки непрерывно выводится 00...0
//
// = Параметры =
// DW [1]: ширина информационной шины i и блоков b(k)
// CW [2]: ширина управляющей шины s и логарифм количества блоков b(k)
module demux(i, s, o);
  parameter DW = 1;
  parameter CW = 2;
  localparam N = 2**CW;
  input [DW-1:0] i;
  input [CW-1:0] s;
  output [DW*N-1:0] o;
  
  reg [DW-1:0] b[0:N-1];
  
  always @(*)
  begin : switch_block
    integer k;
    for(k = 0; k < N; k = k + 1)
      b[k] = {{DW{1'b0}}}; //DW раз повторяй 0
    b[s] = i;
  end
  
  genvar k;
  for(k = 0; k < N; k = k + 1)
    assign o[DW*(N-k)-1:DW*(N-1-k)] = b[k];
endmodule
